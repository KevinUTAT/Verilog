`timescale 1ns / 1ns 

module Lab2p3(SW, HEX0);
	input [3:0] SW;
	output [6:0] HEX0;
	
	hexDecoder hd0(
				.C(SW),
				.H(HEX0)
				);
endmodule			


	
module hexDecoder(C, H);
	input [3:0] C;
	output [6:0] H;
	
	//assigning value to each light
	assign H[0] = (C[3] | C[2] | C[1] | ~C[0]) & (C[3] | ~C[2] | C[1] | C[0]) &
		(~C[3] | C[2] | ~C[1] | ~C[0]) & (~C[3] | ~C[2] | ~C[1] | C[0]);
		
	assign H[1] = (C[3] | ~C[2] | C[1] | ~C[0]) & (C[3] | ~C[2] | ~C[1] | C[0]) & 
		(~C[3] | C[2] | ~C[1] | ~C[0]) & (~C[3] | ~C[2] | C[1] | C[0]) & 
		(~C[3] | ~C[2] | ~C[1] | C[0]) & (~C[3] | ~C[2] | ~C[1] | ~C[0]);
		
	assign H[2] = (C[3] | C[2] | ~C[1] | C[0]) & (~C[3] | ~C[2] | C[1] | C[0]) & 
		(~C[3] | ~C[2] | ~C[1] | C[0]) & (~C[3] | ~C[2] | ~C[1] | ~C[0]);
		
	assign H[3] = (C[3] | C[2] | C[1] | ~C[0]) & (C[3] | ~C[2] | C[1] | C[0]) & 
		(C[3] | ~C[2] | ~C[1] | ~C[0]) & (~C[3] | C[2] | C[1] | ~C[0]) & 
		(~C[3] | C[2] | ~C[1] | C[0]) & (~C[3] | ~C[2] | ~C[1] | ~C[0]);
		
	assign H[4] = (C[3] | C[2] | C[1] | ~C[0]) & (C[3] | C[2] | ~C[1] | ~C[0]) & 
		(C[3] | ~C[2] | C[1] | C[0]) & (C[3] | ~C[2] | C[1] | ~C[0]) & 
		(C[3] | ~C[2] | ~C[1] | ~C[0]) & (~C[3] | C[2] | C[1] | ~C[0]);
		
	assign H[5] = (C[3] | C[2] | C[1] | ~C[0]) & (C[3] | C[2] | ~C[1] | C[0]) & 
		(C[3] | C[2] | ~C[1] | ~C[0]) & (C[3] | ~C[2] | ~C[1] | ~C[0]) & 
		(~C[3] | ~C[2] | C[1] | ~C[0]);
		
	assign H[6] = (C[3] | C[2] | C[1] | C[0]) & (C[3] | C[2] | C[1] | ~C[0]) & 
		(C[3] | ~C[2] | ~C[1] | ~C[0]) & (~C[3] | ~C[2] | C[1] | C[0]);
		
endmodule
